library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD_UNSIGNED.all;  

entity imem is
 port
 (
  pc:   in  STD_LOGIC_VECTOR(31 downto 0);
  inst: out STD_LOGIC_VECTOR(31 downto 0)
 );
end;

architecture Behavioral of imem is
 type Instruction is array (0 to 15) of std_logic_vector(31 downto 0);
 constant rom_data: Instruction:=(
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000",
"00100001001010000000000000100000"
 );
begin
 process is
 begin
  loop
   inst <= rom_data(to_integer(pc)/4);
   wait on pc;
  end loop;
 end process;
end;