library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD_UNSIGNED.all;  

entity imem is
 port
 (
  pc:   in  STD_LOGIC_VECTOR(31 downto 0);
  inst: out STD_LOGIC_VECTOR(31 downto 0)
 );
end;

architecture Behavioral of imem is
 type Instruction is array (0 to 31) of std_logic_vector(31 downto 0);
 constant rom_data: Instruction:=(
  "10000000000000000000000000000000",
  "01000000000000000000000000000000",
  "00100000000000000000000000000000",
  "00010000000000000000000000000000",
  "00001000000000000000000000000000",
  "00000100000000000000000000000000",
  "00000010000000000000000000000000",
  "00000001000000000000000000000000",
  "00000000100000000000000000000000",
  "00000000010000000000000000000000",
  "00000000001000000000000000000000",
  "00000000000100000000000000000000",
  "00000000000010000000000000000000",
  "00000000000001000000000000000000",
  "00000000000000100000000000000000",
  "00000000000000010000000000000000",
  "00000000000000001000000000000000",
  "00000000000000000100000000000000",
  "00000000000000000010000000000000",
  "00000000000000000001000000000000",
  "00000000000000000000100000000000",
  "00000000000000000000010000000000",
  "00000000000000000000001000000000",
  "00000000000000000000000100000000",
  "00000000000000000000000010000000",
  "00000000000000000000000001000000",
  "00000000000000000000000000100000",
  "00000000000000000000000000010000",
  "00000000000000000000000000001000",
  "00000000000000000000000000000100",
  "00000000000000000000000000000010",
  "00000000000000000000000000000001"
 );
begin
 process is
 begin
  loop
   inst <= rom_data(to_integer(pc)/4);
   wait on pc;
  end loop;
 end process;
end;